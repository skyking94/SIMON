////////////////////////////////////////////////////////////////////////////////////////////////////
//
//			RIGHT SHIFT MODULE - PARAMETERIZED
//
////////////////////////////////////////////////////////////////////////////////////////////////////

module right_shifter #(parameter WORD_SIZE=64, SHIFT_COUNT=1)
		(
		input		[WORD_SIZE-1:0]		data_in,
		output		[WORD_SIZE-1:0]		data_out
		);


//--------------------------------------------------------------------------------------------------
//					Assignment Operations
//--------------------------------------------------------------------------------------------------
	
assign data_out = data_in >> SHIFT_COUNT;


endmodule // right_shifter