////////////////////////////////////////////////////////////////////////////////////////////////////
//
//			LEFT SHIFT MODULE - PARAMETERIZED
//
////////////////////////////////////////////////////////////////////////////////////////////////////

module left_shifter #(parameter BLOCK_SIZE=64, SHIFT_COUNT=1)
		(
		input			[BLOCK_SIZE-1:0]			data_in,
		output			[BLOCK_SIZE-1:0]			data_out
		);

//--------------------------------------------------------------------------------------------------
//					Assignment Operations
//--------------------------------------------------------------------------------------------------
assign data_count = data_in << SHIFT_COUNT;



endmodule
